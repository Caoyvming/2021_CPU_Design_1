module mux16_2to1_tb();

//Generate Inputs
reg       [15:0]       D_IN0;
reg       [15:0]       D_IN1;
reg       [15:0]       D_IN2;
reg       [15:0]       D_IN3;
reg       [1:0]          SEL;

//Capture Outputs
wire      [15:0]       D_OUT;

// Instantiate the Unit Under Test (UUT)
mux16_4to1 uut(
    .SEL    (SEL),
    .D_IN0  (D_IN0),
    .D_IN1  (D_IN1),
    .D_IN2  (D_IN2),
    .D_IN3  (D_IN3),
    .D_OUT  (D_OUT)
);

//Encourage
initial begin
        // Initialize Inputs
        D_IN0 = 16'b0000000000000000;
        D_IN1 = 16'b0000000000000000;
        D_IN2 = 16'b0000000000000000;
        D_IN3 = 16'b0000000000000000;
        SEL   = 2'b00               ;

        // Wait 100 ns for global reset to finish
        #100;
        // Add stimulus here
        D_IN0 <= 16'b0000000000000001;
        D_IN1 <= 16'b1000000000000000;
        D_IN2 <= 16'b0000000000000001;
        D_IN3 <= 16'b1000000000000000;
        SEL   = 2'b00                ;

        #100;
        D_IN0 <= 16'b0000000000000010;
        D_IN1 <= 16'b0100000000000000;
        D_IN2 <= 16'b0000000000000010;
        D_IN3 <= 16'b0100000000000000;
        SEL   = 2'b01                ;

        #100;
        D_IN0 <= 16'b0000000000000100;
        D_IN1 <= 16'b0010000000000000;
        D_IN2 <= 16'b0000000000000100;
        D_IN3 <= 16'b0010000000000000;
        SEL   = 2'b10                ;

        #100;
        D_IN0 <= 16'b0000000000001000;
        D_IN1 <= 16'b0001000000000000;
        D_IN2 <= 16'b0000000000001000;
        D_IN3 <= 16'b0001000000000000;
        SEL   = 2'b11                ;
 
        #100;
        D_IN0 <= 16'b0000000000010000;
        D_IN1 <= 16'b0000100000000000;
        D_IN2 <= 16'b0000000000010000;
        D_IN3 <= 16'b0000100000000000;
        SEL   = 2'b00                ;
 
        #100;
        D_IN0 <= 16'b0000000000100000;
        D_IN1 <= 16'b0000010000000000;
        D_IN2 <= 16'b0000000000100000;
        D_IN3 <= 16'b0000010000000000;
        SEL   = 2'b01                ;

        #100;
        D_IN0 <= 16'b0000000001000000;
        D_IN1 <= 16'b0000001000000000;
        D_IN2 <= 16'b0000000001000000;
        D_IN3 <= 16'b0000001000000000;
        SEL   = 2'b10                ;

        #100;
        D_IN0 <= 16'b0000000010000000;
        D_IN1 <= 16'b0000000100000000;
        D_IN2 <= 16'b0000000010000000;
        D_IN3 <= 16'b0000000100000000;
        SEL   = 2'b11                ;
    end
endmodule